module subbytes(
    input [127:0]in_state,
    output [127:0]out_state
);
endmodule