module key_expansion(
    input clk,
    input rst_n,
    input start,
    input [3:0]round,
    input [127:0]key_in,
    output [127:0]round_key
);
endmodule