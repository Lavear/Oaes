module aes_datapath(
    input clk, 
    input rst_n,
    input final_round,
    input [127:0]round_key,
    input [127:0]state_in,
    output [127:0]state_out
);
endmodule