module state_reg(
    input clk,
    input rst_n,
    input enable,
    input [127:0]next_state,
    output reg [127:0]state
);
endmodule